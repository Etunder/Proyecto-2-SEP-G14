library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FFT_tb is
-- Testbench entities do not have ports.
end entity FFT_tb;

architecture tb of FFT_tb is
    -- Component Declaration for the FFT module
    component FFT
        Port (
            clk             : in  std_logic;
            rst             : in  std_logic;
            start           : in std_logic;
            sample_vector   : in  std_logic_vector(2047 downto 0);
            fft_output      : out std_logic_vector(383 downto 0);
            fft_processing_done : out std_logic;
            ROM_data        : in  std_logic_vector(63 downto 0);
            addr            : out std_logic_vector(9 downto 0);
            out_state : out std_logic_vector(2 downto 0);
            coef_received_out : out std_logic;
            partial_done_count_out : out std_logic_vector(4 downto 0)
        );
    end component;

    -- Signals for Interconnecting the Testbench and the FFT
    signal tb_clk   : std_logic := '0';
    signal tb_rst   : std_logic := '0';
    signal tb_sample_vector : std_logic_vector(2047 downto 0) := (others => '0');
    signal tb_fft_output    : std_logic_vector(383 downto 0);
    signal tb_fft_processing_done : std_logic;
    signal tb_ROM_data  : std_logic_vector(63 downto 0);
    signal tb_addr      : std_logic_vector(9 downto 0);
    signal tb_start     : std_logic := '0';
    signal tb_state     : std_logic_vector(2 downto 0);
    signal tb_coef      : std_logic;
    signal tb_partial_done_count : std_logic_vector(4 downto 0);
   
    -- Clock period definition
    constant clk_period : time := 10 ns;
begin
    -- Instantiate the Module Under Test (MUT)
    uut: FFT
        port map (
            clk => tb_clk,
            rst => tb_rst,
            start => tb_start,
            sample_vector => tb_sample_vector,
            fft_output => tb_fft_output,
            fft_processing_done => tb_fft_processing_done,
            ROM_data => tb_ROM_data,
            addr => tb_addr,
            out_state => tb_state, 
            coef_received_out => tb_coef,
            partial_done_count_out => tb_partial_done_count
        );

    -- Clock process
    clk_process : process
    begin
        tb_clk <= '0';
        wait for clk_period/2;
        tb_clk <= '1';
        wait for clk_period/2;
    end process;

    -- Reset process
    rst_process : process
    begin
        tb_start <= '0';
        wait for 20 ns;
        tb_start <= '1';
        wait for 20 ns;
        tb_start <= '0';
        wait;
    end process;

    -- Simulated ROM process
    rom_process : process(tb_addr)
    begin
        -- Define your ROM data based on the address
        case tb_addr is
       when "0000000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0000000001" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0000000010" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0000000011" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0000000100" =>  tb_ROM_data <= "1010010101010011110010011100101010111111100000000000000000000000";
       when "0000000101" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0000000110" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0000000111" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0000001000" =>  tb_ROM_data <= "1011111110000000000000000000000000100101110100111100100111001010";
       when "0000001001" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0000001010" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0000001011" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0000001100" =>  tb_ROM_data <= "0010011000011110110101110101100000111111100000000000000000000000";
       when "0000001101" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0000001110" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0000001111" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0000010000" =>  tb_ROM_data <= "0011111110000000000000000000000010100110010100111100100111001010";
       when "0000010001" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0000010010" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0000010011" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0000010100" =>  tb_ROM_data <= "1010011101000010001011110000111110111111100000000000000000000000";
       when "0000010101" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0000010110" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0000010111" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0000011000" =>  tb_ROM_data <= "1011111110000000000000000000000000100110100111101101011101011000";
       when "0000011001" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0000011010" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0000011011" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0000011100" =>  tb_ROM_data <= "1010011000001101010111101101111000111111100000000000000000000000";
       when "0000011101" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0000011110" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0000011111" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0000100000" =>  tb_ROM_data <= "0011111110000000000000000000000010100110110100111100100111001010";
       when "0000100001" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0000100010" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0000100011" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0000100100" =>  tb_ROM_data <= "1010011101110111001000011000001010111111100000000000000000000000";
       when "0000100101" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0000100110" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0000100111" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0000101000" =>  tb_ROM_data <= "1011111110000000000000000000000000100111110000100010111100001111";
       when "0000101001" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0000101010" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0000101011" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0000101100" =>  tb_ROM_data <= "0010100000000100011001101010111100111111100000000000000000000000";
       when "0000101101" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0000101110" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0000101111" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0000110000" =>  tb_ROM_data <= "0011111110000000000000000000000010100111000111101101011101011000";
       when "0000110001" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0000110010" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0000110011" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0000110100" =>  tb_ROM_data <= "0010011101010011111011000000110010111111100000000000000000000000";
       when "0000110101" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0000110110" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0000110111" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0000111000" =>  tb_ROM_data <= "1011111110000000000000000000000010100110100011010101111011011110";
       when "0000111001" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0000111010" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0000111011" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0000111100" =>  tb_ROM_data <= "0010100010001000110100011010011000111111100000000000000000000000";
       when "0000111101" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0000111110" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0000111111" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0001000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0001000001" =>  tb_ROM_data <= "0011111010010100101000000011000100111111011101001111101000001011";
       when "0001000010" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0001000011" =>  tb_ROM_data <= "1011111101000101111001000000001110111111001000100110011110011001";
       when "0001000100" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0001000101" =>  tb_ROM_data <= "0011111101111110110001000110110100111101110010001011110100110110";
       when "0001000110" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0001000111" =>  tb_ROM_data <= "1011111101100001110001011001100000111110111100010101101011101010";
       when "0001001000" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0001001001" =>  tb_ROM_data <= "0011111011110001010110101110101010111111011000011100010110011000";
       when "0001001010" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0001001011" =>  tb_ROM_data <= "0011110111001000101111010011011000111111011111101100010001101101";
       when "0001001100" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0001001101" =>  tb_ROM_data <= "1011111100100010011001111001100110111111010001011110010000000011";
       when "0001001110" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0001001111" =>  tb_ROM_data <= "0011111101110100111110100000101100111110100101001010000000110001";
       when "0001010000" =>  tb_ROM_data <= "1010011010001101010010000000100000111111100000000000000000000000";
       when "0001010001" =>  tb_ROM_data <= "1011111101110100111110100000101100111110100101001010000000110001";
       when "0001010010" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0001010011" =>  tb_ROM_data <= "0011111100100010011001111001100110111111010001011110010000000011";
       when "0001010100" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0001010101" =>  tb_ROM_data <= "1011110111001000101111010011011000111111011111101100010001101101";
       when "0001010110" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0001010111" =>  tb_ROM_data <= "1011111011110001010110101110101010111111011000011100010110011000";
       when "0001011000" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0001011001" =>  tb_ROM_data <= "0011111101100001110001011001100000111110111100010101101011101010";
       when "0001011010" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0001011011" =>  tb_ROM_data <= "1011111101111110110001000110110100111101110010001011110100110110";
       when "0001011100" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0001011101" =>  tb_ROM_data <= "0011111101000101111001000000001110111111001000100110011110011001";
       when "0001011110" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0001011111" =>  tb_ROM_data <= "1011111010010100101000000011000100111111011101001111101000001011";
       when "0001100000" =>  tb_ROM_data <= "1011111110000000000000000000000010100111000011010100100000001000";
       when "0001100001" =>  tb_ROM_data <= "1011111010010100101000000011000110111111011101001111101000001011";
       when "0001100010" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0001100011" =>  tb_ROM_data <= "0011111101000101111001000000001100111111001000100110011110011001";
       when "0001100100" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0001100101" =>  tb_ROM_data <= "1011111101111110110001000110110110111101110010001011110100110110";
       when "0001100110" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0001100111" =>  tb_ROM_data <= "0011111101100001110001011001100010111110111100010101101011101010";
       when "0001101000" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0001101001" =>  tb_ROM_data <= "1011111011110001010110101110101000111111011000011100010110011000";
       when "0001101010" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0001101011" =>  tb_ROM_data <= "1011110111001000101111010011011010111111011111101100010001101101";
       when "0001101100" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0001101101" =>  tb_ROM_data <= "0011111100100010011001111001100100111111010001011110010000000011";
       when "0001101110" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0001101111" =>  tb_ROM_data <= "1011111101110100111110100000101110111110100101001010000000110001";
       when "0001110000" =>  tb_ROM_data <= "1010011110010110000010011111101010111111100000000000000000000000";
       when "0001110001" =>  tb_ROM_data <= "0011111101110100111110100000101110111110100101001010000000110001";
       when "0001110010" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0001110011" =>  tb_ROM_data <= "1011111100100010011001111001100100111111010001011110010000000011";
       when "0001110100" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0001110101" =>  tb_ROM_data <= "0011110111001000101111010011011010111111011111101100010001101101";
       when "0001110110" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0001110111" =>  tb_ROM_data <= "0011111011110001010110101110101000111111011000011100010110011000";
       when "0001111000" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0001111001" =>  tb_ROM_data <= "1011111101100001110001011001100010111110111100010101101011101010";
       when "0001111010" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0001111011" =>  tb_ROM_data <= "0011111101111110110001000110110110111101110010001011110100110110";
       when "0001111100" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0001111101" =>  tb_ROM_data <= "1011111101000101111001000000001100111111001000100110011110011001";
       when "0001111110" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0001111111" =>  tb_ROM_data <= "0011111010010100101000000011000110111111011101001111101000001011";
       when "0010000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0010000001" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0010000010" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0010000011" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0010000100" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0010000101" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0010000110" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0010000111" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0010001000" =>  tb_ROM_data <= "1010010111110111000101100001011110111111100000000000000000000000";
       when "0010001001" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0010001010" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0010001011" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0010001100" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0010001101" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0010001110" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0010001111" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0010010000" =>  tb_ROM_data <= "1011111110000000000000000000000000100110011101110001011000010111";
       when "0010010001" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0010010010" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0010010011" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0010010100" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0010010101" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0010010110" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0010010111" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0010011000" =>  tb_ROM_data <= "1010011000001101010111101101111000111111100000000000000000000000";
       when "0010011001" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0010011010" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0010011011" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0010011100" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0010011101" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0010011110" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0010011111" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0010100000" =>  tb_ROM_data <= "0011111110000000000000000000000010100110111101110001011000010111";
       when "0010100001" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0010100010" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0010100011" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0010100100" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0010100101" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0010100110" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0010100111" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0010101000" =>  tb_ROM_data <= "1010011110001101001101101110011110111111100000000000000000000000";
       when "0010101001" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0010101010" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0010101011" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0010101100" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0010101101" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0010101110" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0010101111" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0010110000" =>  tb_ROM_data <= "1011111110000000000000000000000010100110100011010101111011011110";
       when "0010110001" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0010110010" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0010110011" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0010110100" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0010110101" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0010110110" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0010110111" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0010111000" =>  tb_ROM_data <= "0010100000010110000011001101010100111111100000000000000000000000";
       when "0010111001" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0010111010" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0010111011" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0010111100" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0010111101" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0010111110" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0010111111" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0011000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0011000001" =>  tb_ROM_data <= "0011110111001000101111010011011000111111011111101100010001101101";
       when "0011000010" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0011000011" =>  tb_ROM_data <= "1011111010010100101000000011000110111111011101001111101000001011";
       when "0011000100" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0011000101" =>  tb_ROM_data <= "0011111011110001010110101110101000111111011000011100010110011000";
       when "0011000110" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0011000111" =>  tb_ROM_data <= "1011111100100010011001111001100110111111010001011110010000000011";
       when "0011001000" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0011001001" =>  tb_ROM_data <= "0011111101000101111001000000001100111111001000100110011110011001";
       when "0011001010" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0011001011" =>  tb_ROM_data <= "1011111101100001110001011001100010111110111100010101101011101010";
       when "0011001100" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0011001101" =>  tb_ROM_data <= "0011111101110100111110100000101100111110100101001010000000110001";
       when "0011001110" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0011001111" =>  tb_ROM_data <= "1011111101111110110001000110110110111101110010001011110100110110";
       when "0011010000" =>  tb_ROM_data <= "1010011101000010001011110000111110111111100000000000000000000000";
       when "0011010001" =>  tb_ROM_data <= "0011111101111110110001000110110110111101110010001011110100110110";
       when "0011010010" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0011010011" =>  tb_ROM_data <= "1011111101110100111110100000101100111110100101001010000000110001";
       when "0011010100" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0011010101" =>  tb_ROM_data <= "0011111101100001110001011001100010111110111100010101101011101010";
       when "0011010110" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0011010111" =>  tb_ROM_data <= "1011111101000101111001000000001100111111001000100110011110011001";
       when "0011011000" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0011011001" =>  tb_ROM_data <= "0011111100100010011001111001100110111111010001011110010000000011";
       when "0011011010" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0011011011" =>  tb_ROM_data <= "1011111011110001010110101110101000111111011000011100010110011000";
       when "0011011100" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0011011101" =>  tb_ROM_data <= "0011111010010100101000000011000110111111011101001111101000001011";
       when "0011011110" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0011011111" =>  tb_ROM_data <= "1011110111001000101111010011011000111111011111101100010001101101";
       when "0011100000" =>  tb_ROM_data <= "1011111110000000000000000000000000100111110000100010111100001111";
       when "0011100001" =>  tb_ROM_data <= "1011110111001000101111010011011010111111011111101100010001101101";
       when "0011100010" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0011100011" =>  tb_ROM_data <= "0011111010010100101000000011000100111111011101001111101000001011";
       when "0011100100" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0011100101" =>  tb_ROM_data <= "1011111011110001010110101110101010111111011000011100010110011000";
       when "0011100110" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0011100111" =>  tb_ROM_data <= "0011111100100010011001111001100100111111010001011110010000000011";
       when "0011101000" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0011101001" =>  tb_ROM_data <= "1011111101000101111001000000001110111111001000100110011110011001";
       when "0011101010" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0011101011" =>  tb_ROM_data <= "0011111101100001110001011001100000111110111100010101101011101010";
       when "0011101100" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0011101101" =>  tb_ROM_data <= "1011111101110100111110100000101110111110100101001010000000110001";
       when "0011101110" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0011101111" =>  tb_ROM_data <= "0011111101111110110001000110110100111101110010001011110100110110";
       when "0011110000" =>  tb_ROM_data <= "0010011010001101000110100101101100111111100000000000000000000000";
       when "0011110001" =>  tb_ROM_data <= "1011111101111110110001000110110100111101110010001011110100110110";
       when "0011110010" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0011110011" =>  tb_ROM_data <= "0011111101110100111110100000101110111110100101001010000000110001";
       when "0011110100" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0011110101" =>  tb_ROM_data <= "1011111101100001110001011001100000111110111100010101101011101010";
       when "0011110110" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0011110111" =>  tb_ROM_data <= "0011111101000101111001000000001110111111001000100110011110011001";
       when "0011111000" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0011111001" =>  tb_ROM_data <= "1011111100100010011001111001100100111111010001011110010000000011";
       when "0011111010" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0011111011" =>  tb_ROM_data <= "0011111011110001010110101110101010111111011000011100010110011000";
       when "0011111100" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0011111101" =>  tb_ROM_data <= "1011111010010100101000000011000100111111011101001111101000001011";
       when "0011111110" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0011111111" =>  tb_ROM_data <= "0011110111001000101111010011011010111111011111101100010001101101";
       when "0100000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0100000001" =>  tb_ROM_data <= "0010010010001101001100010011001000111111100000000000000000000000";
       when "0100000010" =>  tb_ROM_data <= "1011111110000000000000000000000000100101000011010011000100110010";
       when "0100000011" =>  tb_ROM_data <= "1010010101010011110010011100101010111111100000000000000000000000";
       when "0100000100" =>  tb_ROM_data <= "0011111110000000000000000000000010100101100011010011000100110010";
       when "0100000101" =>  tb_ROM_data <= "0010010110110000011111010111111000111111100000000000000000000000";
       when "0100000110" =>  tb_ROM_data <= "1011111110000000000000000000000000100101110100111100100111001010";
       when "0100000111" =>  tb_ROM_data <= "1010010111110111000101100001011110111111100000000000000000000000";
       when "0100001000" =>  tb_ROM_data <= "0011111110000000000000000000000010100110000011010011000100110010";
       when "0100001001" =>  tb_ROM_data <= "0010011000011110110101110101100000111111100000000000000000000000";
       when "0100001010" =>  tb_ROM_data <= "1011111110000000000000000000000000100110001100000111110101111110";
       when "0100001011" =>  tb_ROM_data <= "1010011100110000100010001110100110111111100000000000000000000000";
       when "0100001100" =>  tb_ROM_data <= "0011111110000000000000000000000010100110010100111100100111001010";
       when "0100001101" =>  tb_ROM_data <= "1010011010001101010010000000100000111111100000000000000000000000";
       when "0100001110" =>  tb_ROM_data <= "1011111110000000000000000000000000100110011101110001011000010111";
       when "0100001111" =>  tb_ROM_data <= "1010011101000010001011110000111110111111100000000000000000000000";
       when "0100010000" =>  tb_ROM_data <= "0011111110000000000000000000000010100110100011010011000100110010";
       when "0100010001" =>  tb_ROM_data <= "1010011001010011111101110111011100111111100000000000000000000000";
       when "0100010010" =>  tb_ROM_data <= "1011111110000000000000000000000000100110100111101101011101011000";
       when "0100010011" =>  tb_ROM_data <= "1010011101010011110101010011010110111111100000000000000000000000";
       when "0100010100" =>  tb_ROM_data <= "0011111110000000000000000000000010100110101100000111110101111110";
       when "0100010101" =>  tb_ROM_data <= "1010011000001101010111101101111000111111100000000000000000000000";
       when "0100010110" =>  tb_ROM_data <= "1011111110000000000000000000000000100111101100001000100011101001";
       when "0100010111" =>  tb_ROM_data <= "1010011101100101011110110101110010111111100000000000000000000000";
       when "0100011000" =>  tb_ROM_data <= "0011111110000000000000000000000010100110110100111100100111001010";
       when "0100011001" =>  tb_ROM_data <= "1010010110001101100011001000101000111111100000000000000000000000";
       when "0100011010" =>  tb_ROM_data <= "1011111110000000000000000000000010100111000011010100100000001000";
       when "0100011011" =>  tb_ROM_data <= "1010011101110111001000011000001010111111100000000000000000000000";
       when "0100011100" =>  tb_ROM_data <= "0011111110000000000000000000000010100110111101110001011000010111";
       when "0100011101" =>  tb_ROM_data <= "1010000100110110101100001101101100111111100000000000000000000000";
       when "0100011110" =>  tb_ROM_data <= "1011111110000000000000000000000000100111110000100010111100001111";
       when "0100011111" =>  tb_ROM_data <= "1010011110000100011000111101010010111111100000000000000000000000";
       when "0100100000" =>  tb_ROM_data <= "0011111110000000000000000000000010100111000011010011000100110010";
       when "0100100001" =>  tb_ROM_data <= "0010010110001100110101011101100100111111100000000000000000000000";
       when "0100100010" =>  tb_ROM_data <= "1011111110000000000000000000000010100110110100111111011101110111";
       when "0100100011" =>  tb_ROM_data <= "1010011110001101001101101110011110111111100000000000000000000000";
       when "0100100100" =>  tb_ROM_data <= "0011111110000000000000000000000010100111000111101101011101011000";
       when "0100100101" =>  tb_ROM_data <= "0010011000001101000000111000010100111111100000000000000000000000";
       when "0100100110" =>  tb_ROM_data <= "1011111110000000000000000000000000100111110100111101010100110101";
       when "0100100111" =>  tb_ROM_data <= "1010011110010110000010011111101010111111100000000000000000000000";
       when "0100101000" =>  tb_ROM_data <= "0011111110000000000000000000000010100111001100000111110101111110";
       when "0100101001" =>  tb_ROM_data <= "0010100000001101001110011100001000111111100000000000000000000000";
       when "0100101010" =>  tb_ROM_data <= "1011111110000000000000000000000010100110100011010101111011011110";
       when "0100101011" =>  tb_ROM_data <= "1010011110011110110111010000110110111111100000000000000000000000";
       when "0100101100" =>  tb_ROM_data <= "0011111110000000000000000000000010101000001100001000100011101001";
       when "0100101101" =>  tb_ROM_data <= "0010011010001101000110100101101100111111100000000000000000000000";
       when "0100101110" =>  tb_ROM_data <= "1011111110000000000000000000000000100111111001010111101101011100";
       when "0100101111" =>  tb_ROM_data <= "0010011100110000100111111011111110111111100000000000000000000000";
       when "0100110000" =>  tb_ROM_data <= "0011111110000000000000000000000010100111010100111100100111001010";
       when "0100110001" =>  tb_ROM_data <= "0010100000010110000011001101010100111111100000000000000000000000";
       when "0100110010" =>  tb_ROM_data <= "1011111110000000000000000000000010100110000011011000110010001010";
       when "0100110011" =>  tb_ROM_data <= "1010011110110000100000110011010010111111100000000000000000000000";
       when "0100110100" =>  tb_ROM_data <= "0011111110000000000000000000000000100111100011010100100000001000";
       when "0100110101" =>  tb_ROM_data <= "0010011011010011101100101111010000111111100000000000000000000000";
       when "0100110110" =>  tb_ROM_data <= "1011111110000000000000000000000000100111111101110010000110000010";
       when "0100110111" =>  tb_ROM_data <= "0010011100001101010100110111001110111111100000000000000000000000";
       when "0100111000" =>  tb_ROM_data <= "0011111110000000000000000000000010100111011101110001011000010111";
       when "0100111001" =>  tb_ROM_data <= "0010100000011110110111111110100000111111100000000000000000000000";
       when "0100111010" =>  tb_ROM_data <= "1011111110000000000000000000000010100001101101101011000011011011";
       when "0100111011" =>  tb_ROM_data <= "1010011111000010001010010101101010111111100000000000000000000000";
       when "0100111100" =>  tb_ROM_data <= "0011111110000000000000000000000010101000010000100010111100001111";
       when "0100111101" =>  tb_ROM_data <= "0010011100001101001001011100011100111111100000000000000000000000";
       when "0100111110" =>  tb_ROM_data <= "1011111110000000000000000000000000101000000001000110001111010100";
       when "0100111111" =>  tb_ROM_data <= "0010011011010100000011100100110110111111100000000000000000000000";
       when "0101000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0101000001" =>  tb_ROM_data <= "1011110111001000101111010011011000111111011111101100010001101101";
       when "0101000010" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0101000011" =>  tb_ROM_data <= "0011111010010100101000000011000110111111011101001111101000001011";
       when "0101000100" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0101000101" =>  tb_ROM_data <= "1011111011110001010110101110101000111111011000011100010110011000";
       when "0101000110" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0101000111" =>  tb_ROM_data <= "0011111100100010011001111001100110111111010001011110010000000011";
       when "0101001000" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0101001001" =>  tb_ROM_data <= "1011111101000101111001000000001100111111001000100110011110011001";
       when "0101001010" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0101001011" =>  tb_ROM_data <= "0011111101100001110001011001100010111110111100010101101011101010";
       when "0101001100" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0101001101" =>  tb_ROM_data <= "1011111101110100111110100000101100111110100101001010000000110001";
       when "0101001110" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0101001111" =>  tb_ROM_data <= "0011111101111110110001000110110110111101110010001011110100110110";
       when "0101010000" =>  tb_ROM_data <= "1010011001010011111101110111011100111111100000000000000000000000";
       when "0101010001" =>  tb_ROM_data <= "1011111101111110110001000110110110111101110010001011110100110110";
       when "0101010010" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0101010011" =>  tb_ROM_data <= "0011111101110100111110100000101100111110100101001010000000110001";
       when "0101010100" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0101010101" =>  tb_ROM_data <= "1011111101100001110001011001100010111110111100010101101011101010";
       when "0101010110" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0101010111" =>  tb_ROM_data <= "0011111101000101111001000000001100111111001000100110011110011001";
       when "0101011000" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0101011001" =>  tb_ROM_data <= "1011111100100010011001111001100110111111010001011110010000000011";
       when "0101011010" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0101011011" =>  tb_ROM_data <= "0011111011110001010110101110101000111111011000011100010110011000";
       when "0101011100" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0101011101" =>  tb_ROM_data <= "1011111010010100101000000011000110111111011101001111101000001011";
       when "0101011110" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0101011111" =>  tb_ROM_data <= "0011110111001000101111010011011000111111011111101100010001101101";
       when "0101100000" =>  tb_ROM_data <= "1011111110000000000000000000000010100110110100111111011101110111";
       when "0101100001" =>  tb_ROM_data <= "0011110111001000101111010011011010111111011111101100010001101101";
       when "0101100010" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0101100011" =>  tb_ROM_data <= "1011111010010100101000000011000100111111011101001111101000001011";
       when "0101100100" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0101100101" =>  tb_ROM_data <= "0011111011110001010110101110101010111111011000011100010110011000";
       when "0101100110" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0101100111" =>  tb_ROM_data <= "1011111100100010011001111001100100111111010001011110010000000011";
       when "0101101000" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0101101001" =>  tb_ROM_data <= "0011111101000101111001000000001110111111001000100110011110011001";
       when "0101101010" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0101101011" =>  tb_ROM_data <= "1011111101100001110001011001100000111110111100010101101011101010";
       when "0101101100" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0101101101" =>  tb_ROM_data <= "0011111101110100111110100000101110111110100101001010000000110001";
       when "0101101110" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0101101111" =>  tb_ROM_data <= "1011111101111110110001000110110100111101110010001011110100110110";
       when "0101110000" =>  tb_ROM_data <= "1010011110110000100000110011010010111111100000000000000000000000";
       when "0101110001" =>  tb_ROM_data <= "0011111101111110110001000110110100111101110010001011110100110110";
       when "0101110010" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0101110011" =>  tb_ROM_data <= "1011111101110100111110100000101110111110100101001010000000110001";
       when "0101110100" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0101110101" =>  tb_ROM_data <= "0011111101100001110001011001100000111110111100010101101011101010";
       when "0101110110" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0101110111" =>  tb_ROM_data <= "1011111101000101111001000000001110111111001000100110011110011001";
       when "0101111000" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0101111001" =>  tb_ROM_data <= "0011111100100010011001111001100100111111010001011110010000000011";
       when "0101111010" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0101111011" =>  tb_ROM_data <= "1011111011110001010110101110101010111111011000011100010110011000";
       when "0101111100" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0101111101" =>  tb_ROM_data <= "0011111010010100101000000011000100111111011101001111101000001011";
       when "0101111110" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0101111111" =>  tb_ROM_data <= "1011110111001000101111010011011010111111011111101100010001101101";
       when "0110000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0110000001" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0110000010" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0110000011" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0110000100" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0110000101" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0110000110" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0110000111" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0110001000" =>  tb_ROM_data <= "0010011000011110110101110101100000111111100000000000000000000000";
       when "0110001001" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0110001010" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0110001011" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0110001100" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0110001101" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0110001110" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0110001111" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0110010000" =>  tb_ROM_data <= "1011111110000000000000000000000000100110100111101101011101011000";
       when "0110010001" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0110010010" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0110010011" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0110010100" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0110010101" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0110010110" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0110010111" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0110011000" =>  tb_ROM_data <= "1010011101110111001000011000001010111111100000000000000000000000";
       when "0110011001" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0110011010" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0110011011" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0110011100" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0110011101" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0110011110" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0110011111" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0110100000" =>  tb_ROM_data <= "0011111110000000000000000000000010100111000111101101011101011000";
       when "0110100001" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0110100010" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0110100011" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0110100100" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0110100101" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0110100110" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0110100111" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0110101000" =>  tb_ROM_data <= "0010011010001101000110100101101100111111100000000000000000000000";
       when "0110101001" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0110101010" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0110101011" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0110101100" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0110101101" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0110101110" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0110101111" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0110110000" =>  tb_ROM_data <= "1011111110000000000000000000000000100111111101110010000110000010";
       when "0110110001" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0110110010" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0110110011" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0110110100" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0110110101" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0110110110" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0110110111" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0110111000" =>  tb_ROM_data <= "0010011011010100000011100100110110111111100000000000000000000000";
       when "0110111001" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0110111010" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0110111011" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0110111100" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0110111101" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0110111110" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0110111111" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0111000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "0111000001" =>  tb_ROM_data <= "1011111010010100101000000011000100111111011101001111101000001011";
       when "0111000010" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "0111000011" =>  tb_ROM_data <= "0011111101000101111001000000001110111111001000100110011110011001";
       when "0111000100" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "0111000101" =>  tb_ROM_data <= "1011111101111110110001000110110100111101110010001011110100110110";
       when "0111000110" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "0111000111" =>  tb_ROM_data <= "0011111101100001110001011001100000111110111100010101101011101010";
       when "0111001000" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "0111001001" =>  tb_ROM_data <= "1011111011110001010110101110101010111111011000011100010110011000";
       when "0111001010" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "0111001011" =>  tb_ROM_data <= "1011110111001000101111010011011000111111011111101100010001101101";
       when "0111001100" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "0111001101" =>  tb_ROM_data <= "0011111100100010011001111001100110111111010001011110010000000011";
       when "0111001110" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "0111001111" =>  tb_ROM_data <= "1011111101110100111110100000101100111110100101001010000000110001";
       when "0111010000" =>  tb_ROM_data <= "1010011101010011110101010011010110111111100000000000000000000000";
       when "0111010001" =>  tb_ROM_data <= "0011111101110100111110100000101100111110100101001010000000110001";
       when "0111010010" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "0111010011" =>  tb_ROM_data <= "1011111100100010011001111001100110111111010001011110010000000011";
       when "0111010100" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "0111010101" =>  tb_ROM_data <= "0011110111001000101111010011011000111111011111101100010001101101";
       when "0111010110" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "0111010111" =>  tb_ROM_data <= "0011111011110001010110101110101010111111011000011100010110011000";
       when "0111011000" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "0111011001" =>  tb_ROM_data <= "1011111101100001110001011001100000111110111100010101101011101010";
       when "0111011010" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "0111011011" =>  tb_ROM_data <= "0011111101111110110001000110110100111101110010001011110100110110";
       when "0111011100" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "0111011101" =>  tb_ROM_data <= "1011111101000101111001000000001110111111001000100110011110011001";
       when "0111011110" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "0111011111" =>  tb_ROM_data <= "0011111010010100101000000011000100111111011101001111101000001011";
       when "0111100000" =>  tb_ROM_data <= "1011111110000000000000000000000000100111110100111101010100110101";
       when "0111100001" =>  tb_ROM_data <= "0011111010010100101000000011000110111111011101001111101000001011";
       when "0111100010" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "0111100011" =>  tb_ROM_data <= "1011111101000101111001000000001100111111001000100110011110011001";
       when "0111100100" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "0111100101" =>  tb_ROM_data <= "0011111101111110110001000110110110111101110010001011110100110110";
       when "0111100110" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "0111100111" =>  tb_ROM_data <= "1011111101100001110001011001100010111110111100010101101011101010";
       when "0111101000" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "0111101001" =>  tb_ROM_data <= "0011111011110001010110101110101000111111011000011100010110011000";
       when "0111101010" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "0111101011" =>  tb_ROM_data <= "0011110111001000101111010011011010111111011111101100010001101101";
       when "0111101100" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "0111101101" =>  tb_ROM_data <= "1011111100100010011001111001100100111111010001011110010000000011";
       when "0111101110" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "0111101111" =>  tb_ROM_data <= "0011111101110100111110100000101110111110100101001010000000110001";
       when "0111110000" =>  tb_ROM_data <= "0010100000011110110111111110100000111111100000000000000000000000";
       when "0111110001" =>  tb_ROM_data <= "1011111101110100111110100000101110111110100101001010000000110001";
       when "0111110010" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "0111110011" =>  tb_ROM_data <= "0011111100100010011001111001100100111111010001011110010000000011";
       when "0111110100" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "0111110101" =>  tb_ROM_data <= "1011110111001000101111010011011010111111011111101100010001101101";
       when "0111110110" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "0111110111" =>  tb_ROM_data <= "1011111011110001010110101110101000111111011000011100010110011000";
       when "0111111000" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "0111111001" =>  tb_ROM_data <= "0011111101100001110001011001100010111110111100010101101011101010";
       when "0111111010" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "0111111011" =>  tb_ROM_data <= "1011111101111110110001000110110110111101110010001011110100110110";
       when "0111111100" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "0111111101" =>  tb_ROM_data <= "0011111101000101111001000000001100111111001000100110011110011001";
       when "0111111110" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "0111111111" =>  tb_ROM_data <= "1011111010010100101000000011000110111111011101001111101000001011";
       when "1000000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "1000000001" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1000000010" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1000000011" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1000000100" =>  tb_ROM_data <= "0010010110110000011111010111111000111111100000000000000000000000";
       when "1000000101" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1000000110" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1000000111" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1000001000" =>  tb_ROM_data <= "1011111110000000000000000000000000100110001100000111110101111110";
       when "1000001001" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1000001010" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1000001011" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1000001100" =>  tb_ROM_data <= "1010011101000010001011110000111110111111100000000000000000000000";
       when "1000001101" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1000001110" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1000001111" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1000010000" =>  tb_ROM_data <= "0011111110000000000000000000000010100110101100000111110101111110";
       when "1000010001" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1000010010" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1000010011" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1000010100" =>  tb_ROM_data <= "1010010110001101100011001000101000111111100000000000000000000000";
       when "1000010101" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1000010110" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1000010111" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1000011000" =>  tb_ROM_data <= "1011111110000000000000000000000000100111110000100010111100001111";
       when "1000011001" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1000011010" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1000011011" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1000011100" =>  tb_ROM_data <= "1010011110001101001101101110011110111111100000000000000000000000";
       when "1000011101" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1000011110" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1000011111" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1000100000" =>  tb_ROM_data <= "0011111110000000000000000000000010100111001100000111110101111110";
       when "1000100001" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1000100010" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1000100011" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1000100100" =>  tb_ROM_data <= "0010011010001101000110100101101100111111100000000000000000000000";
       when "1000100101" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1000100110" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1000100111" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1000101000" =>  tb_ROM_data <= "1011111110000000000000000000000010100110000011011000110010001010";
       when "1000101001" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1000101010" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1000101011" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1000101100" =>  tb_ROM_data <= "1010100001011100101010110010001110111111100000000000000000000000";
       when "1000101101" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1000101110" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1000101111" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1000110000" =>  tb_ROM_data <= "0011111110000000000000000000000010101000010000100010111100001111";
       when "1000110001" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1000110010" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1000110011" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1000110100" =>  tb_ROM_data <= "1010011110110000100110100000101000111111100000000000000000000000";
       when "1000110101" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1000110110" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1000110111" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1000111000" =>  tb_ROM_data <= "1011111110000000000000000000000000101000000011010011011011100111";
       when "1000111001" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1000111010" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1000111011" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1000111100" =>  tb_ROM_data <= "1010011111100101011101011010011010111111100000000000000000000000";
       when "1000111101" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1000111110" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1000111111" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1001000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "1001000001" =>  tb_ROM_data <= "1011111011110001010110101110101000111111011000011100010110011000";
       when "1001000010" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "1001000011" =>  tb_ROM_data <= "0011111101111110110001000110110110111101110010001011110100110110";
       when "1001000100" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1001000101" =>  tb_ROM_data <= "1011111100100010011001111001100110111111010001011110010000000011";
       when "1001000110" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "1001000111" =>  tb_ROM_data <= "1011111010010100101000000011000100111111011101001111101000001011";
       when "1001001000" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1001001001" =>  tb_ROM_data <= "0011111101110100111110100000101110111110100101001010000000110001";
       when "1001001010" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "1001001011" =>  tb_ROM_data <= "1011111101000101111001000000001110111111001000100110011110011001";
       when "1001001100" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1001001101" =>  tb_ROM_data <= "1011110111001000101111010011011000111111011111101100010001101101";
       when "1001001110" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "1001001111" =>  tb_ROM_data <= "0011111101100001110001011001100010111110111100010101101011101010";
       when "1001010000" =>  tb_ROM_data <= "1010011000001101010111101101111000111111100000000000000000000000";
       when "1001010001" =>  tb_ROM_data <= "1011111101100001110001011001100010111110111100010101101011101010";
       when "1001010010" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "1001010011" =>  tb_ROM_data <= "0011110111001000101111010011011000111111011111101100010001101101";
       when "1001010100" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1001010101" =>  tb_ROM_data <= "0011111101000101111001000000001110111111001000100110011110011001";
       when "1001010110" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "1001010111" =>  tb_ROM_data <= "1011111101110100111110100000101110111110100101001010000000110001";
       when "1001011000" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1001011001" =>  tb_ROM_data <= "0011111010010100101000000011000100111111011101001111101000001011";
       when "1001011010" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "1001011011" =>  tb_ROM_data <= "0011111100100010011001111001100110111111010001011110010000000011";
       when "1001011100" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1001011101" =>  tb_ROM_data <= "1011111101111110110001000110110110111101110010001011110100110110";
       when "1001011110" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "1001011111" =>  tb_ROM_data <= "0011111011110001010110101110101000111111011000011100010110011000";
       when "1001100000" =>  tb_ROM_data <= "1011111110000000000000000000000010100110100011010101111011011110";
       when "1001100001" =>  tb_ROM_data <= "0011111011110001010110101110101010111111011000011100010110011000";
       when "1001100010" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "1001100011" =>  tb_ROM_data <= "1011111101111110110001000110110100111101110010001011110100110110";
       when "1001100100" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1001100101" =>  tb_ROM_data <= "0011111100100010011001111001100100111111010001011110010000000011";
       when "1001100110" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "1001100111" =>  tb_ROM_data <= "0011111010010100101000000011000110111111011101001111101000001011";
       when "1001101000" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1001101001" =>  tb_ROM_data <= "1011111101110100111110100000101100111110100101001010000000110001";
       when "1001101010" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "1001101011" =>  tb_ROM_data <= "0011111101000101111001000000001100111111001000100110011110011001";
       when "1001101100" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1001101101" =>  tb_ROM_data <= "0011110111001000101111010011011010111111011111101100010001101101";
       when "1001101110" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "1001101111" =>  tb_ROM_data <= "1011111101100001110001011001100000111110111100010101101011101010";
       when "1001110000" =>  tb_ROM_data <= "0010011011010100000011100100110110111111100000000000000000000000";
       when "1001110001" =>  tb_ROM_data <= "0011111101100001110001011001100000111110111100010101101011101010";
       when "1001110010" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "1001110011" =>  tb_ROM_data <= "1011110111001000101111010011011010111111011111101100010001101101";
       when "1001110100" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1001110101" =>  tb_ROM_data <= "1011111101000101111001000000001100111111001000100110011110011001";
       when "1001110110" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "1001110111" =>  tb_ROM_data <= "0011111101110100111110100000101100111110100101001010000000110001";
       when "1001111000" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1001111001" =>  tb_ROM_data <= "1011111010010100101000000011000110111111011101001111101000001011";
       when "1001111010" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "1001111011" =>  tb_ROM_data <= "1011111100100010011001111001100100111111010001011110010000000011";
       when "1001111100" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1001111101" =>  tb_ROM_data <= "0011111101111110110001000110110100111101110010001011110100110110";
       when "1001111110" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "1001111111" =>  tb_ROM_data <= "1011111011110001010110101110101010111111011000011100010110011000";
       when "1010000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "1010000001" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "1010000010" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1010000011" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "1010000100" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1010000101" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "1010000110" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1010000111" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "1010001000" =>  tb_ROM_data <= "1010011100110000100010001110100110111111100000000000000000000000";
       when "1010001001" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "1010001010" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1010001011" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "1010001100" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1010001101" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "1010001110" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1010001111" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "1010010000" =>  tb_ROM_data <= "1011111110000000000000000000000000100111101100001000100011101001";
       when "1010010001" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "1010010010" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1010010011" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "1010010100" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1010010101" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "1010010110" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1010010111" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "1010011000" =>  tb_ROM_data <= "0010010110001100110101011101100100111111100000000000000000000000";
       when "1010011001" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "1010011010" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1010011011" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "1010011100" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1010011101" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "1010011110" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1010011111" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "1010100000" =>  tb_ROM_data <= "0011111110000000000000000000000010101000001100001000100011101001";
       when "1010100001" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "1010100010" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1010100011" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "1010100100" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1010100101" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "1010100110" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1010100111" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "1010101000" =>  tb_ROM_data <= "0010011100001101010100110111001110111111100000000000000000000000";
       when "1010101001" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "1010101010" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1010101011" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "1010101100" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1010101101" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "1010101110" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1010101111" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "1010110000" =>  tb_ROM_data <= "1011111110000000000000000000000000100110000011001101010111011001";
       when "1010110001" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "1010110010" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1010110011" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "1010110100" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1010110101" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "1010110110" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1010110111" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "1010111000" =>  tb_ROM_data <= "0010011101010011101111100101111100111111100000000000000000000000";
       when "1010111001" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "1010111010" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1010111011" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "1010111100" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1010111101" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "1010111110" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1010111111" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "1011000000" =>  tb_ROM_data <= "0011111110000000000000000000000000000000000000000000000000000000";
       when "1011000001" =>  tb_ROM_data <= "1011111100100010011001111001100100111111010001011110010000000011";
       when "1011000010" =>  tb_ROM_data <= "1011111001000111110001011100001010111111011110110001010010111110";
       when "1011000011" =>  tb_ROM_data <= "0011111101100001110001011001100000111110111100010101101011101010";
       when "1011000100" =>  tb_ROM_data <= "1011111101101100100000110101111000111110110000111110111100010101";
       when "1011000101" =>  tb_ROM_data <= "0011111010010100101000000011000110111111011101001111101000001011";
       when "1011000110" =>  tb_ROM_data <= "0011111100001110001110011101101000111111010101001101101100110001";
       when "1011000111" =>  tb_ROM_data <= "1011111101111110110001000110110110111101110010001011110100110110";
       when "1011001000" =>  tb_ROM_data <= "0011111100110101000001001111001110111111001101010000010011110011";
       when "1011001001" =>  tb_ROM_data <= "0011110111001000101111010011011000111111011111101100010001101101";
       when "1011001010" =>  tb_ROM_data <= "1011111101010100110110110011000110111111000011100011100111011010";
       when "1011001011" =>  tb_ROM_data <= "0011111101110100111110100000101110111110100101001010000000110001";
       when "1011001100" =>  tb_ROM_data <= "1011111011000011111011110001010100111111011011001000001101011110";
       when "1011001101" =>  tb_ROM_data <= "1011111011110001010110101110101010111111011000011100010110011000";
       when "1011001110" =>  tb_ROM_data <= "0011111101111011000101001011111000111110010001111100010111000010";
       when "1011001111" =>  tb_ROM_data <= "1011111101000101111001000000001100111111001000100110011110011001";
       when "1011010000" =>  tb_ROM_data <= "1010011101100101011110110101110010111111100000000000000000000000";
       when "1011010001" =>  tb_ROM_data <= "0011111101000101111001000000001100111111001000100110011110011001";
       when "1011010010" =>  tb_ROM_data <= "1011111101111011000101001011111000111110010001111100010111000010";
       when "1011010011" =>  tb_ROM_data <= "0011111011110001010110101110101010111111011000011100010110011000";
       when "1011010100" =>  tb_ROM_data <= "0011111011000011111011110001010100111111011011001000001101011110";
       when "1011010101" =>  tb_ROM_data <= "1011111101110100111110100000101110111110100101001010000000110001";
       when "1011010110" =>  tb_ROM_data <= "0011111101010100110110110011000110111111000011100011100111011010";
       when "1011010111" =>  tb_ROM_data <= "1011110111001000101111010011011000111111011111101100010001101101";
       when "1011011000" =>  tb_ROM_data <= "1011111100110101000001001111001110111111001101010000010011110011";
       when "1011011001" =>  tb_ROM_data <= "0011111101111110110001000110110110111101110010001011110100110110";
       when "1011011010" =>  tb_ROM_data <= "1011111100001110001110011101101000111111010101001101101100110001";
       when "1011011011" =>  tb_ROM_data <= "1011111010010100101000000011000110111111011101001111101000001011";
       when "1011011100" =>  tb_ROM_data <= "0011111101101100100000110101111000111110110000111110111100010101";
       when "1011011101" =>  tb_ROM_data <= "1011111101100001110001011001100000111110111100010101101011101010";
       when "1011011110" =>  tb_ROM_data <= "0011111001000111110001011100001010111111011110110001010010111110";
       when "1011011111" =>  tb_ROM_data <= "0011111100100010011001111001100100111111010001011110010000000011";
       when "1011100000" =>  tb_ROM_data <= "1011111110000000000000000000000000100111111001010111101101011100";
       when "1011100001" =>  tb_ROM_data <= "0011111100100010011001111001100110111111010001011110010000000011";
       when "1011100010" =>  tb_ROM_data <= "0011111001000111110001011100001000111111011110110001010010111110";
       when "1011100011" =>  tb_ROM_data <= "1011111101100001110001011001100010111110111100010101101011101010";
       when "1011100100" =>  tb_ROM_data <= "0011111101101100100000110101111010111110110000111110111100010101";
       when "1011100101" =>  tb_ROM_data <= "1011111010010100101000000011000100111111011101001111101000001011";
       when "1011100110" =>  tb_ROM_data <= "1011111100001110001110011101101010111111010101001101101100110001";
       when "1011100111" =>  tb_ROM_data <= "0011111101111110110001000110110100111101110010001011110100110110";
       when "1011101000" =>  tb_ROM_data <= "1011111100110101000001001111001100111111001101010000010011110011";
       when "1011101001" =>  tb_ROM_data <= "1011110111001000101111010011011010111111011111101100010001101101";
       when "1011101010" =>  tb_ROM_data <= "0011111101010100110110110011000100111111000011100011100111011010";
       when "1011101011" =>  tb_ROM_data <= "1011111101110100111110100000101100111110100101001010000000110001";
       when "1011101100" =>  tb_ROM_data <= "0011111011000011111011110001010110111111011011001000001101011110";
       when "1011101101" =>  tb_ROM_data <= "0011111011110001010110101110101000111111011000011100010110011000";
       when "1011101110" =>  tb_ROM_data <= "1011111101111011000101001011111010111110010001111100010111000010";
       when "1011101111" =>  tb_ROM_data <= "0011111101000101111001000000001110111111001000100110011110011001";
       when "1011110000" =>  tb_ROM_data <= "0010011100110000011100100001001100111111100000000000000000000000";
       when "1011110001" =>  tb_ROM_data <= "1011111101000101111001000000001110111111001000100110011110011001";
       when "1011110010" =>  tb_ROM_data <= "0011111101111011000101001011111010111110010001111100010111000010";
       when "1011110011" =>  tb_ROM_data <= "1011111011110001010110101110101000111111011000011100010110011000";
       when "1011110100" =>  tb_ROM_data <= "1011111011000011111011110001010110111111011011001000001101011110";
       when "1011110101" =>  tb_ROM_data <= "0011111101110100111110100000101100111110100101001010000000110001";
       when "1011110110" =>  tb_ROM_data <= "1011111101010100110110110011000100111111000011100011100111011010";
       when "1011110111" =>  tb_ROM_data <= "0011110111001000101111010011011010111111011111101100010001101101";
       when "1011111000" =>  tb_ROM_data <= "0011111100110101000001001111001100111111001101010000010011110011";
       when "1011111001" =>  tb_ROM_data <= "1011111101111110110001000110110100111101110010001011110100110110";
       when "1011111010" =>  tb_ROM_data <= "0011111100001110001110011101101010111111010101001101101100110001";
       when "1011111011" =>  tb_ROM_data <= "0011111010010100101000000011000100111111011101001111101000001011";
       when "1011111100" =>  tb_ROM_data <= "1011111101101100100000110101111010111110110000111110111100010101";
       when "1011111101" =>  tb_ROM_data <= "0011111101100001110001011001100010111110111100010101101011101010";
       when "1011111110" =>  tb_ROM_data <= "1011111001000111110001011100001000111111011110110001010010111110";
       when "1011111111" =>  tb_ROM_data <= "1011111100100010011001111001100110111111010001011110010000000011";
       when others => tb_ROM_data <= (others => '0');
        end case;
    end process;

    -- Test stimulus process
    stim_proc: process
    begin
        -- Initialize Inputs
        tb_sample_vector (31 downto 0) <= "01000000010000000000000000000000";

        -- Wait for global reset to finish
        wait for 50 ns;
        

        -- Insert stimulus here, e.g., setting sample_vector values

        wait;
    end process;

end architecture tb;
